Graph := G (1, 1, 1)